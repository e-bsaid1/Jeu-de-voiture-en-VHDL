library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--Une procédure est un type de sous-programme en VHDL qui peut nous aider à éviter la répétition du code. 
--Il est parfois nécessaire d'effectuer des opérations identiques à plusieurs endroits de la conception.


PACKAGE DELIMITATIONS_TRONCONS IS
PROCEDURE DELIMITATIONS_TRONCON
(
  SIGNAL DELIMITATIONS_TRONCON_current_pos_X,DELIMITATIONS_TRONCON_current_pos_Y,Xpos,Ypos:IN INTEGER;
  SIGNAL RGB_DELIMITATIONS_TRONCON:OUT STD_LOGIC_VECTOR(3 downto 0);
  SIGNAL DRAWING_DELIMITATIONS_TRONCON: OUT STD_LOGIC;
  CONSTANT LARGEUR_DELIMITATIONS_TRONCON:INTEGER;
  CONSTANT LONGUEUR_DELIMITATIONS_TRONCON:INTEGER
  );
END DELIMITATIONS_TRONCONS;



PACKAGE BODY DELIMITATIONS_TRONCONS IS
PROCEDURE DELIMITATIONS_TRONCON
(
  SIGNAL DELIMITATIONS_TRONCON_current_pos_X,DELIMITATIONS_TRONCON_current_pos_Y,Xpos,Ypos:IN INTEGER;
  SIGNAL RGB_DELIMITATIONS_TRONCON:OUT STD_LOGIC_VECTOR(3 downto 0);
  SIGNAL DRAWING_DELIMITATIONS_TRONCON: OUT STD_LOGIC;
  CONSTANT LARGEUR_DELIMITATIONS_TRONCON:INTEGER;
  CONSTANT LONGUEUR_DELIMITATIONS_TRONCON:INTEGER)
  IS
  
---------- Si le compteur atteint se situe dans les X et Y mentionnés ci-dessous, faire apparaitre le gazon
  BEGIN
    IF((DELIMITATIONS_TRONCON_current_pos_X>Xpos) AND (DELIMITATIONS_TRONCON_current_pos_X<(Xpos+LARGEUR_DELIMITATIONS_TRONCON)) AND (DELIMITATIONS_TRONCON_current_pos_Y>Ypos) AND (DELIMITATIONS_TRONCON_current_pos_Y<(Ypos+LONGUEUR_DELIMITATIONS_TRONCON)))THEN
	    RGB_DELIMITATIONS_TRONCON<="1111";
	    DRAWING_DELIMITATIONS_TRONCON<='1';
		 
		 ELSE 
		 DRAWING_DELIMITATIONS_TRONCON<='0';
 END IF;
 
END DELIMITATIONS_TRONCON;
END DELIMITATIONS_TRONCONS;